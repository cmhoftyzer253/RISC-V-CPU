import cpu_consts::*;

module multiply (
    input logic [63:0] opr_a_i,
    input logic [63:0] opr_b_i,

    input logic [2:0] mult_func_i,

    output logic [63:0] mult_res_o
);

    logic [63:0] mult_res_o;

endmodule