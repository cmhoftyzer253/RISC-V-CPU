module branch_control (

);



endmodule;