import cpu_consts::*;

module divide (
    input logic [63:0] opr_a_i,
    input logic [63:0] opr_b_i,

    input logic [2:0] div_func_i,

    output logic [63:0] div_res_o
);

    output logic [63:0] div_res_o;

endmodule